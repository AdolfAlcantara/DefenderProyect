/* verilator lint_off WIDTH */
module MemDecoder (
    input [31:0] virtAddr, //! Virtual address
    output [12:0] physAddr, //! Physical address
    output invalidAddr //! Invalid address
);

endmodule
