`define ADDI   6'h08
`define ADDIU  6'h09
`define ANDI   6'h0C
`define ORI    6'h0D
`define LUI    6'h0F
`define ADD    6'h20
`define ADDU   6'h21
`define SUB    6'h22
`define SUBU   6'h23
`define AND    6'h24
`define OR     6'h25
`define SLT    6'h2A
`define SLTI   6'h0A
`define SLTU   6'h2B
`define SLTIU  6'h0B
`define LW     6'h23
`define SW     6'h2B
`define BEQ    6'h04
`define BNE    6'h05
`define JUMP   6'h02
`define XOR    6'h26
`define XORI   6'h0E

`define LH     6'h21
`define LHU    6'h25
`define LB     6'h20
`define LBU    6'h24
`define SH     6'h29
`define SB     6'h28
