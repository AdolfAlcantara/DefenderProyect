/* verilator lint_off WIDTH */
/* verilator lint_off UNUSED */
module PCDecoder (
    input [31:0] virtPC, //! Virtual PC
    output [11:0] physPC, //! Physical PC
    output invalidPC // Invalid program counter
);

endmodule
